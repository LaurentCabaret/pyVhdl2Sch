hello world in the new file
and another line
